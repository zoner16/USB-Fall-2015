sumanamugothu@Sumans-MacBook-Pro.local.10605